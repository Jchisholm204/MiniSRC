// ALU Verilog Header File

// Control Parameters
`define CTRL_ALU_ADD 4'h0
`define CTRL_ALU_SUB 4'h1
`define CTRL_ALU_OR  4'h2
`define CTRL_ALU_XOR 4'h3
`define CTRL_ALU_AND 4'h4
`define CTRL_ALU_MUL 4'h5
`define CTRL_ALU_DIV 4'h6
`define CTRL_ALU_SLL 4'h7
`define CTRL_ALU_SRL 4'h8
`define CTRL_ALU_SRA 4'h9
`define CTRL_ALU_ROR 4'hA
`define CTRL_ALU_ROL 4'hB
