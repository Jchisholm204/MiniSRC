/**
* Jacob Chisholm
* DE2 VGA Parameters
*   Designed for a 640x480 resolution signal
*/

`define VGA_WIDTH 32'd640
`define VGA_WIDTH 32'd640
