`ifndef _constants_vh_
`define _constants_vh_

`define START_PC_ADDRESS 32'h00000000

`endif