module ControlUnit(
    
);

endmodule