module miniSRC();

Processor proc(

)

endmodule