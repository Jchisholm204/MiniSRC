`ifndef _constants_vh_
`define _constants_vh_

`define START_PC_ADDRESS 32'h00000000
// Set to 1 for simulation (makes life easier)
// Must be set to 4 
`define PC_INCREMENT 32'h00000004

`endif
